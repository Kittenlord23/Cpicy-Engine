default -> type_setting_vsync[True] -> type_setting_frame_delay[60] -> layers[1] -> type_text[] -> type_rect[[288,173,173,231,255,255,255,1,00000001,1,0]::[670,309,197,319,255,255,255,1,00000005,1,0]::] -> type_line[] -> type_image[] -> type_rect_wall[[287,171,176,234,1,00000002]::[1,1083,1914,148,0,00000003]::[671,307,195,318,1,00000006]::] -> end <->