default -> type_setting_vsync[True] -> type_setting_frame_delay[60] -> layers[1] -> type_text[] -> type_rect[[878,465,264,209,184,0,253,0,00000009,1,0]::] -> type_line[] -> type_image[[167,405,403,201,0,1,SPACESHIP_1.png,00000002,1,0]::] -> type_rect_wall[[171,515,324,82,1,00000003]::[-202,1,202,1084,0,00000004]::[-2,1079,1926,137,0,00000005]::[1921,-3,159,1083,0,00000006]::[-12,-118,1930,115,0,00000007]::[990,-285,1,8,0,00000008]::[874,461,270,216,0,000000010]::] -> end <->